# ====================================================================
#
#      hal_arm_arm9_ep93xx.cdl
#
#      Cirrus Logic ARM9/EP93XX platform HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#                                                                          
# -------------------------------------------                              
# The contents of this file are subject to the Red Hat eCos Public License 
# Version 1.1 (the "License"); you may not use this file except in         
# compliance with the License.  You may obtain a copy of the License at    
# http://www.redhat.com/                                                   
#                                                                          
# Software distributed under the License is distributed on an "AS IS"      
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the 
# License for the specific language governing rights and limitations under 
# the License.                                                             
#                                                                          
# The Original Code is eCos - Embedded Configurable Operating System,      
# released September 30, 1998.                                             
#                                                                          
# The Initial Developer of the Original Code is Red Hat.                   
# Portions created by Red Hat are                                          
# Copyright (C) 1998, 1999, 2000, 2001 Red Hat, Inc.                             
# All Rights Reserved.                                                     
# -------------------------------------------                              
#                                                                          
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Original data:  gthomas
# Contributors:   paul.jordan
# Date:           2001-04-11
#
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_HAL_ARM_ARM9_EP93XX {
    display       "Cirrus Logic ARM9/EP93xx evaluation board"
    parent        CYGPKG_HAL_ARM_ARM9
    requires      CYGPKG_HAL_ARM_ARM9_ARM920T
    hardware
    include_dir   cyg/hal
    define_header hal_arm_arm9_ep93xx.h
    description   "This HAL platform package provides generic
        support for the Cirrus Logic EP93xx based boards."

    compile       ep93xx_misc.c hal_diag.c terk.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_arm_arm9.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_arm9_ep93xx.h>"
        puts $::cdl_header "#define HAL_PLATFORM_CPU    \"ARM920T\""
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        default_value {"RAM"}
        legal_values  {"RAM" "ROMRAM" }
        no_define
        define -file system.h CYG_HAL_STARTUP
        description   "
           When targetting the EP93xx eval board it is possible to build
           the system for either RAM bootstrap or ROM bootstrap(s). Select
           'ram' when building programs to load into RAM using eCos GDB
           stubs.  Select 'rom' when building a stand-alone application
           which will be put into ROM, or for the special case of
           building the eCos GDB stubs themselves."
    }

    cdl_option CYGHWR_HAL_ARM_EDB93XX_VARIANT {
        display       "Cirrus Logic processor variant"
        flavor        data
        legal_values  { "EP9301" "EP9302" "EP9307" "EP9312" "EP9315" "EP9315A"}
        default_value { "EP9312" }
        description   "
            The Cirrus Logic processor variant."
        define -file system.h CYGHWR_HAL_ARM_EDB93XX_VARIANT
    }

    cdl_option CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT {
        display       "Cirrus Logic board variant"
        flavor        data
        legal_values  { "EDB9301" "EDB9302" "EDB9307" "EDB9312" "EDB9315" "EDB9315A"}
        default_value { CYGHWR_HAL_ARM_EDB93XX_VARIANT == "EP9301" ? "EDB9301" : \
                        CYGHWR_HAL_ARM_EDB93XX_VARIANT == "EP9302" ? "EDB9302" : \
                        CYGHWR_HAL_ARM_EDB93XX_VARIANT == "EP9307" ? "EDB9307" : \
                        CYGHWR_HAL_ARM_EDB93XX_VARIANT == "EP9312" ? "EDB9312" : \
                        CYGHWR_HAL_ARM_EDB93XX_VARIANT == "EP9315" ? "EDB9315" : \
                        CYGHWR_HAL_ARM_EDB93XX_VARIANT == "EP9315A" ? "EDB9315A" : \
                        "" }
        description   "
            The board type which uses a Cirrus Logic processor variant."
        define -file system.h CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT
	    
        define_proc {
            puts $::cdl_header ""
            puts $::cdl_header "#ifdef CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT_EDB9301"
            puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Cirrus Logic EDB9301 Board\""
            puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"Rev A\""
            puts $::cdl_header "#define HAL_PLATFORM_EP9301"
            puts $::cdl_header "#define HAL_PLATFORM_MACHINE_TYPE  462"
            puts $::cdl_header "#define CYGHWR_REDBOOT_ARM_TRAMPOLINE_ADDRESS 0x00001f00"
            puts $::cdl_header "#endif //CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT_EDB9301"
            puts $::cdl_header ""
            puts $::cdl_header "#ifdef CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT_EDB9302"
            puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Cirrus Logic EDB9302 Board\""
            puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"Rev A\""
            puts $::cdl_header "#define HAL_PLATFORM_EP9302"
            puts $::cdl_header "#define HAL_PLATFORM_MACHINE_TYPE  538"
            puts $::cdl_header "#define CYGHWR_REDBOOT_ARM_TRAMPOLINE_ADDRESS 0x00001f00"
            puts $::cdl_header "#endif //CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT_EDB9302"
            puts $::cdl_header ""
            puts $::cdl_header "#ifdef CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT_EDB9307"
            puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Cirrus Logic EDB9307 Board\""
            puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"Rev A\""
            puts $::cdl_header "#define HAL_PLATFORM_EP9307"
            puts $::cdl_header "#define HAL_PLATFORM_MACHINE_TYPE  607"
            puts $::cdl_header "#define CYGHWR_REDBOOT_ARM_TRAMPOLINE_ADDRESS 0x00001f00"
            puts $::cdl_header "#endif //CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT_EDB9307"
            puts $::cdl_header ""
            puts $::cdl_header "#ifdef CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT_EDB9312"
            puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Cirrus Logic EDB9312 Board\""
            puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"Rev A\""
            puts $::cdl_header "#define HAL_PLATFORM_EP9312"
            puts $::cdl_header "#define HAL_PLATFORM_MACHINE_TYPE  451"
            puts $::cdl_header "#define CYGHWR_REDBOOT_ARM_TRAMPOLINE_ADDRESS 0x00001f00"
            puts $::cdl_header "#endif //CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT_EDB9312"
            puts $::cdl_header ""
            puts $::cdl_header "#ifdef CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT_EDB9315"
            puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Cirrus Logic EDB9315 Board\""
            puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"Rev A\""
            puts $::cdl_header "#define HAL_PLATFORM_EP9315"
            puts $::cdl_header "#define HAL_PLATFORM_MACHINE_TYPE  463"
            puts $::cdl_header "#define CYGHWR_REDBOOT_ARM_TRAMPOLINE_ADDRESS 0x00001f00"
            puts $::cdl_header "#endif //CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT_EDB9315"
            puts $::cdl_header ""
            puts $::cdl_header "#ifdef CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT_EDB9315A"
            puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"Cirrus Logic EDB9315A Board\""
            puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"Rev A\""
            puts $::cdl_header "#define HAL_PLATFORM_EP9315"
            puts $::cdl_header "#define HAL_PLATFORM_MACHINE_TYPE  772"
            puts $::cdl_header "#define CYGHWR_REDBOOT_ARM_TRAMPOLINE_ADDRESS 0x00001f00"
            puts $::cdl_header "#endif //CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT_EDB9315A"
            puts $::cdl_header ""
	    }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { 
          CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9301" ? 
            (CYG_HAL_STARTUP == "RAM" ? "arm_arm9_edb9301_ram" : \
             CYG_HAL_STARTUP == "ROMRAM" ? "arm_arm9_edb9301_romram" : "BOGUS.mlt" ) : \
          CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9302" ? 
            (CYG_HAL_STARTUP == "RAM" ? "arm_arm9_edb9302_ram" : \
             CYG_HAL_STARTUP == "ROMRAM" ? "arm_arm9_edb9302_romram" : "BOGUS.mlt" ) : \
          CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9307" ? 
            (CYG_HAL_STARTUP == "RAM" ? "arm_arm9_edb9307_ram" : \
             CYG_HAL_STARTUP == "ROMRAM" ? "arm_arm9_edb9307_romram" : "BOGUS.mlt" ) : \
          CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9312" ? 
            (CYG_HAL_STARTUP == "RAM" ? "arm_arm9_edb9312_ram" : \
             CYG_HAL_STARTUP == "ROMRAM" ? "arm_arm9_edb9312_romram" : "BOGUS.mlt" ) : \
          CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9315" ? 
            (CYG_HAL_STARTUP == "RAM" ? "arm_arm9_edb9315_ram" : \
             CYG_HAL_STARTUP == "ROMRAM" ? "arm_arm9_edb9315_romram" : "BOGUS.mlt" ) : \
          CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9315A" ? 
            (CYG_HAL_STARTUP == "RAM" ? "arm_arm9_edb9315a_ram" : \
             CYG_HAL_STARTUP == "ROMRAM" ? "arm_arm9_edb9315a_romram" : "BOGUS.mlt" ) : \
          "BOGUS.mlt"
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { 
              CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9301" ?
                (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_edb9301_ram.ldi>" :  \
                 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_arm9_edb9301_romram.ldi>" :  "BOGUS.ldi" ) : \
              CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9302" ?
                (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_edb9302_ram.ldi>" :  \
                 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_arm9_edb9302_romram.ldi>" :  "BOGUS.ldi" ) : \
              CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9307" ?
                (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_edb9307_ram.ldi>" :  \
                 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_arm9_edb9307_romram.ldi>" :  "BOGUS.ldi" ) : \
              CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9312" ?
                (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_edb9312_ram.ldi>" :  \
                 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_arm9_edb9312_romram.ldi>" :  "BOGUS.ldi" ) : \
              CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9315" ?
                (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_edb9315_ram.ldi>" :  \
                 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_arm9_edb9315_romram.ldi>" :  "BOGUS.ldi" ) : \
              CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9315A" ?
                (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_edb9315a_ram.ldi>" :  \
                 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_arm9_edb9315a_romram.ldi>" :  "BOGUS.ldi" ) : \
              "BOGUS.ldi" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated {
              CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9301" ?
                (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_edb9301_ram.h>" :  \
                 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_arm9_edb9301_romram.h>" :  "BOGUS.h" ) : \
              CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9302" ?
                (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_edb9302_ram.h>" :  \
                 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_arm9_edb9302_romram.h>" :  "BOGUS.h" ) : \
              CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9307" ?
                (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_edb9307_ram.h>" :  \
                 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_arm9_edb9307_romram.h>" :  "BOGUS.h" ) : \
              CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9312" ?
                (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_edb9312_ram.h>" :  \
                 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_arm9_edb9312_romram.h>" :  "BOGUS.h" ) : \
              CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9315" ?
                (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_edb9315_ram.h>" :  \
                 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_arm9_edb9315_romram.h>" :  "BOGUS.h" ) : \
              CYGHWR_HAL_ARM_EDB93XX_BOARD_VARIANT == "EDB9315A" ?
                (CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_arm9_edb9315a_ram.h>" :  \
                 CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_arm_arm9_edb9315a_romram.h>" :  "BOGUS.h" ) : \
              "BOGUS.h" }
        }
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
        no_define

        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    (5120)                    ;# Assumes 512KHz clock
        }
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 57600
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 57600
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   1
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The ep93xx board has three serial ports. This option
            chooses which port will be used to connect to a host
            running GDB."
     }

     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    0
         description      "
            The ep93xx board has three serial ports.  This option
            chooses which port will be used for diagnostic output."
     }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT {
        display      "Default console channel."
        flavor       data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        calculated   0
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        no_define
        description   "
        Global build options including control over
        compiler flags, linker flags and choice of toolchain."

        parent  CYGPKG_NONE

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-Wl,--gc-sections -Wl,-static -g -O2 -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROMRAM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.srec : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) --remove-section=.fixed_vectors $< gdb_module.tmp
                $(OBJCOPY) -O srec --change-address 0x10000000 gdb_module.tmp $@
            }
        }
    }

    cdl_option CYG_HAL_ARM_ARM9_EP93XX_PREAMBLE {
        display       "Include module preamble"
        flavor        bool
        default_value { CYGPKG_REDBOOT && (CYG_HAL_STARTUP == "ROMRAM") }
        description   "
            Enable this option to have the Cirrus Logic format module
            header prepended to the image.  This is required of programs,
            such as RedBoot, which are to be placed in Flash, or for
            those programs which are downloaded using the hardware based
            serial download process."
    }

    cdl_option CYG_HAL_ARM_ARM9_EP93XX_SDRAM_CS {
        display       "Chip select used for SDRAM"
        flavor        data
        legal_values  { "SDCSn0" "SDCSn1" "SDCSn2" "SDCSn3" }
        default_value { CYGHWR_HAL_ARM_EDB93XX_VARIANT == "EP9301" ? "SDCSn3" : \
                        CYGHWR_HAL_ARM_EDB93XX_VARIANT == "EP9302" ? "SDCSn3" : \
                        CYGHWR_HAL_ARM_EDB93XX_VARIANT == "EP9307" ? "SDCSn3" : \
                        CYGHWR_HAL_ARM_EDB93XX_VARIANT == "EP9312" ? "SDCSn3" : \
                        CYGHWR_HAL_ARM_EDB93XX_VARIANT == "EP9315" ? "SDCSn3" : \
                        CYGHWR_HAL_ARM_EDB93XX_VARIANT == "EP9315A" ? "SDCSn0" : \
                        "" }
        description   "
            The SDRAM controller chip select to which the board's SDRAM is
            connected."
        define -file system.h CYG_HAL_ARM_ARM9_EP93XX_SDRAM_CS
    }

    cdl_component CYGPKG_HAL_ARM_ARM9_EP93XX_OPTIONS {
        display "ARM9/EP93XX build options"
        flavor  none
        no_define
        description   "
        Package specific build options including control over
        compiler flags used only in building this package,
        and details of which tests are built."


        cdl_option CYGPKG_HAL_ARM_ARM9_EP93XX_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the ARM9 EP93XX HAL. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_HAL_ARM_ARM9_EP93XX_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the ARM9 EP93XX HAL. These flags are removed from
                the set of global flags if present."
        }

        cdl_option CYGPKG_HAL_ARM_ARM9_EP93XX_TESTS {
            display "ARM9/EP93XX tests"
            flavor  data
            no_define
            calculated { "" }
            description   "
                This option specifies the set of tests for the ARM9 EP93xx HAL."
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires { CYG_HAL_STARTUP == "ROMRAM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "Generic" "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             Firstly there is \"Generic\" support which prevents the HAL
             from overriding the hardware vectors that it does not use, to
             instead allow an installed ROM monitor to handle them. This is
             the most basic support which is likely to be common to most
             implementations of ROM monitor.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
     }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to the various relocated SREC images needed
                         for flash updating."

            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf <PREFIX>/bin/image_hdr.o
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img)
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

}
